`include "myCPU.h"
module MEM_stage(

    );

endmodule
