`include"myCPU.h"
module WB_stage(
	
    );
	
endmodule